module slave_port_tb;

endmodule