module demo();
endmodule