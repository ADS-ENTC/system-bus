module slave_port();

endmodule