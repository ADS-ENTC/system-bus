module master_port_tb;
    
endmodule