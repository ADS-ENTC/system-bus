module master_port (
    
);
    
endmodule